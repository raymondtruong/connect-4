// megafunction wizard: %RAM: 1-PORT%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: altsyncram 

// ============================================================
// File Name: ramTP.v
// Megafunction Name(s):
// 			altsyncram
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 17.0.0 Build 595 04/25/2017 SJ Lite Edition
// ************************************************************


//Copyright (C) 2017  Intel Corporation. All rights reserved.
//Your use of Intel Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Intel Program License 
//Subscription Agreement, the Intel Quartus Prime License Agreement,
//the Intel MegaCore Function License Agreement, or other 
//applicable license agreement, including, without limitation, 
//that your use is for the sole purpose of programming logic 
//devices manufactured by Intel and sold by Intel or its 
//authorized distributors.  Please refer to the applicable 
//agreement for further details.

module GameBoard(Clk, SW, enable);
input Clk;
input enable;
input [9:0] SW;
//input reset_n;
reg [5:0] address = 6'd0;
wire [1:0] out;
reg [98:0] gameBoardSequence = 98'd1;

// Assign registers which will be used to evaluate the current state of the rows in the game board.
wire [13:0] row_0;
wire [13:0] row_1;
wire [13:0] row_2;
wire [13:0] row_3;
wire [13:0] row_4;
wire [13:0] row_5;
wire [13:0] row_6;

assign row_0 = gameBoardSequence[13:0];
assign row_1 = gameBoardSequence[27:14];
assign row_2 = gameBoardSequence[41:28];
assign row_3 = gameBoardSequence[55:42];
assign row_4 = gameBoardSequence[69:56];
assign row_5 = gameBoardSequence[83:70];
assign row_6 = gameBoardSequence[98:84]; 

// Assign registers which will be used to evaluate the current state of the columns in the game board.
wire [13:0] column_0;
wire [13:0] column_1;
wire [13:0] column_2;
wire [13:0] column_3;
wire [13:0] column_4;
wire [13:0] column_5;
wire [13:0] column_6;

assign column_0 = {gameBoardSequence[0], gameBoardSequence[7], gameBoardSequence[14], gameBoardSequence[21], gameBoardSequence[28], gameBoardSequence[35], gameBoardSequence[42]};
assign column_1 = {gameBoardSequence[1], gameBoardSequence[8], gameBoardSequence[15], gameBoardSequence[22], gameBoardSequence[29], gameBoardSequence[36], gameBoardSequence[43]};
assign column_2 = {gameBoardSequence[2], gameBoardSequence[9], gameBoardSequence[16], gameBoardSequence[23], gameBoardSequence[30], gameBoardSequence[37], gameBoardSequence[44]};
assign column_3 = {gameBoardSequence[3], gameBoardSequence[10], gameBoardSequence[17], gameBoardSequence[24], gameBoardSequence[31], gameBoardSequence[38], gameBoardSequence[45]};
assign column_4 = {gameBoardSequence[4], gameBoardSequence[11], gameBoardSequence[18], gameBoardSequence[25], gameBoardSequence[32], gameBoardSequence[39], gameBoardSequence[46]};
assign column_5 = {gameBoardSequence[5], gameBoardSequence[12], gameBoardSequence[19], gameBoardSequence[26], gameBoardSequence[33], gameBoardSequence[40], gameBoardSequence[47]};
assign column_6 = {gameBoardSequence[6], gameBoardSequence[13], gameBoardSequence[20], gameBoardSequence[27], gameBoardSequence[34], gameBoardSequence[41], gameBoardSequence[48]};

// we have (49 * 2) - 24 possible positions and we have 13 2'b00 buffers so we need (74 + 26) = 100 bits
wire [99:0] diagonals;
assign diagonals = {gameBoardSequence[3], gameBoardSequence[11], gameBoardSequence[19], gameBoardSequence[27], 2'b00,  gameBoardSequence[2], 
					gameBoardSequence[10], gameBoardSequence[18], gameBoardSequence[26], gameBoardSequence[34], 2'b00, gameBoardSequence[1], 
					gameBoardSequence[9], gameBoardSequence[17], gameBoardSequence[25], gameBoardSequence[33], gameBoardSequence[41],
					2'b00, gameBoardSequence[0], gameBoardSequence[8], gameBoardSequence[16], gameBoardSequence[24],gameBoardSequence[32], 
					gameBoardSequence[40], gameBoardSequence[48],2'b00, gameBoardSequence[7], gameBoardSequence[15], gameBoardSequence[23],
					gameBoardSequence[31], gameBoardSequence[39], gameBoardSequence[47], 2'b00, gameBoardSequence[14], gameBoardSequence[22], 
					gameBoardSequence[30], gameBoardSequence[38], gameBoardSequence[46], 2'b00, gameBoardSequence[21], gameBoardSequence[29], 
					gameBoardSequence[37], gameBoardSequence[45], 2'b00, gameBoardSequence[21], gameBoardSequence[15], gameBoardSequence[9], 
					gameBoardSequence[3] , 2'b00, gameBoardSequence[28], gameBoardSequence[22], gameBoardSequence[16], gameBoardSequence[10], 
					gameBoardSequence[4], 2'b00, gameBoardSequence[35], gameBoardSequence[29], gameBoardSequence[23], gameBoardSequence[17],
					gameBoardSequence[11], gameBoardSequence[5], 2'b00, gameBoardSequence[42], gameBoardSequence[36], gameBoardSequence[30], 
					gameBoardSequence[24], gameBoardSequence[18], gameBoardSequence[12], gameBoardSequence[6], 2'b00, gameBoardSequence[43], 
					gameBoardSequence[37], gameBoardSequence[31], gameBoardSequence[25], gameBoardSequence[19], gameBoardSequence[13], 2'b00,
					gameBoardSequence[44], gameBoardSequence[38], gameBoardSequence[32], gameBoardSequence[26], gameBoardSequence[20], 2'b00,
					gameBoardSequence[45], gameBoardSequence[39], gameBoardSequence[33], gameBoardSequence[27]};

// Wire which contains all winning combinations 
// we need 100 bits for diagonals, 14 * 14 for the rows and columns and 2 * 14 bit for the buffers = 324 bits
wire [323:0] winningCombinations = {row_0, 2'b00, row_1, 2'b00, row_2, 2'b00, row_3, 2'b00, row_4, 2'b00, row_5, 2'b00, row_6,
								2'b00, column_0, 2'b00, column_1, 2'b00, column_2, 2'b00, column_3, 2'b00, column_4, 2'b00, column_5, 2'b00, column_6,
								2'b00, diagonals};

ramTP ram(
.address(address),
.clock(Clk),
.data(SW[1:0]),
.wren(SW[9]),
.q(out[1:0])
);

// Changes the address synchornously with the clock and resets if the max value is reached or if reset_n is high.
always @(posedge Clk)
begin 
	if (address == 6'd49 || SW[8])
		address <= 6'd0;
	else if (enable)
		gameBoardSequence <= gameBoardSequence << 3;
		gameBoardSequence <= {gameBoardSequence[95:0], out, 1'b0};
		address <= address + 1'd1;
	
end 

endmodule


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module ramTP (
	address,
	clock,
	data,
	wren,
	q);

	input	[5:0]  address;
	input	  clock;
	input	[1:0]  data;
	input	  wren;
	output	[1:0]  q;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
	tri1	  clock;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

	wire [1:0] sub_wire0;
	wire [1:0] q = sub_wire0[1:0];

	altsyncram	altsyncram_component (
				.address_a (address),
				.clock0 (clock),
				.data_a (data),
				.wren_a (wren),
				.q_a (sub_wire0),
				.aclr0 (1'b0),
				.aclr1 (1'b0),
				.address_b (1'b1),
				.addressstall_a (1'b0),
				.addressstall_b (1'b0),
				.byteena_a (1'b1),
				.byteena_b (1'b1),
				.clock1 (1'b1),
				.clocken0 (1'b1),
				.clocken1 (1'b1),
				.clocken2 (1'b1),
				.clocken3 (1'b1),
				.data_b (1'b1),
				.eccstatus (),
				.q_b (),
				.rden_a (1'b1),
				.rden_b (1'b1),
				.wren_b (1'b0));
	defparam
		altsyncram_component.clock_enable_input_a = "BYPASS",
		altsyncram_component.clock_enable_output_a = "BYPASS",
		altsyncram_component.intended_device_family = "Cyclone V",
		altsyncram_component.lpm_hint = "enable_RUNTIME_MOD=NO",
		altsyncram_component.lpm_type = "altsyncram",
		altsyncram_component.numwords_a = 64,
		altsyncram_component.operation_mode = "SINGLE_PORT",
		altsyncram_component.outdata_aclr_a = "NONE",
		altsyncram_component.outdata_reg_a = "UNREGISTERED",
		altsyncram_component.power_up_uninitialized = "FALSE",
		altsyncram_component.read_during_write_mode_port_a = "NEW_DATA_NO_NBE_READ",
		altsyncram_component.widthad_a = 6,
		altsyncram_component.width_a = 2,
		altsyncram_component.width_byteena_a = 1;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: ADDRESSSTALL_A NUMERIC "0"
// Retrieval info: PRIVATE: AclrAddr NUMERIC "0"
// Retrieval info: PRIVATE: AclrByte NUMERIC "0"
// Retrieval info: PRIVATE: AclrData NUMERIC "0"
// Retrieval info: PRIVATE: AclrOutput NUMERIC "0"
// Retrieval info: PRIVATE: BYTE_enable NUMERIC "0"
// Retrieval info: PRIVATE: BYTE_SIZE NUMERIC "8"
// Retrieval info: PRIVATE: BlankMemory NUMERIC "1"
// Retrieval info: PRIVATE: CLOCK_enable_INPUT_A NUMERIC "0"
// Retrieval info: PRIVATE: CLOCK_enable_OUTPUT_A NUMERIC "0"
// Retrieval info: PRIVATE: Clken NUMERIC "0"
// Retrieval info: PRIVATE: DataBusSeparated NUMERIC "1"
// Retrieval info: PRIVATE: IMPLEMENT_IN_LES NUMERIC "0"
// Retrieval info: PRIVATE: INIT_FILE_LAYOUT STRING "PORT_A"
// Retrieval info: PRIVATE: INIT_TO_SIM_X NUMERIC "0"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
// Retrieval info: PRIVATE: JTAG_enableD NUMERIC "0"
// Retrieval info: PRIVATE: JTAG_ID STRING "NONE"
// Retrieval info: PRIVATE: MAXIMUM_DEPTH NUMERIC "0"
// Retrieval info: PRIVATE: MIFfilename STRING ""
// Retrieval info: PRIVATE: NUMWORDS_A NUMERIC "64"
// Retrieval info: PRIVATE: RAM_BLOCK_TYPE NUMERIC "0"
// Retrieval info: PRIVATE: READ_DURING_WRITE_MODE_PORT_A NUMERIC "3"
// Retrieval info: PRIVATE: RegAddr NUMERIC "1"
// Retrieval info: PRIVATE: RegData NUMERIC "1"
// Retrieval info: PRIVATE: RegOutput NUMERIC "0"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: SingleClock NUMERIC "1"
// Retrieval info: PRIVATE: UseDQRAM NUMERIC "1"
// Retrieval info: PRIVATE: WRCONTROL_ACLR_A NUMERIC "0"
// Retrieval info: PRIVATE: WidthAddr NUMERIC "6"
// Retrieval info: PRIVATE: WidthData NUMERIC "2"
// Retrieval info: PRIVATE: rden NUMERIC "0"
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: CONSTANT: CLOCK_enable_INPUT_A STRING "BYPASS"
// Retrieval info: CONSTANT: CLOCK_enable_OUTPUT_A STRING "BYPASS"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
// Retrieval info: CONSTANT: LPM_HINT STRING "enable_RUNTIME_MOD=NO"
// Retrieval info: CONSTANT: LPM_TYPE STRING "altsyncram"
// Retrieval info: CONSTANT: NUMWORDS_A NUMERIC "64"
// Retrieval info: CONSTANT: OPERATION_MODE STRING "SINGLE_PORT"
// Retrieval info: CONSTANT: OUTDATA_ACLR_A STRING "NONE"
// Retrieval info: CONSTANT: OUTDATA_REG_A STRING "UNREGISTERED"
// Retrieval info: CONSTANT: POWER_UP_UNINITIALIZED STRING "FALSE"
// Retrieval info: CONSTANT: READ_DURING_WRITE_MODE_PORT_A STRING "NEW_DATA_NO_NBE_READ"
// Retrieval info: CONSTANT: WIDTHAD_A NUMERIC "6"
// Retrieval info: CONSTANT: WIDTH_A NUMERIC "2"
// Retrieval info: CONSTANT: WIDTH_BYTEENA_A NUMERIC "1"
// Retrieval info: USED_PORT: address 0 0 6 0 INPUT NODEFVAL "address[5..0]"
// Retrieval info: USED_PORT: clock 0 0 0 0 INPUT VCC "clock"
// Retrieval info: USED_PORT: data 0 0 2 0 INPUT NODEFVAL "data[1..0]"
// Retrieval info: USED_PORT: q 0 0 2 0 OUTPUT NODEFVAL "q[1..0]"
// Retrieval info: USED_PORT: wren 0 0 0 0 INPUT NODEFVAL "wren"
// Retrieval info: CONNECT: @address_a 0 0 6 0 address 0 0 6 0
// Retrieval info: CONNECT: @clock0 0 0 0 0 clock 0 0 0 0
// Retrieval info: CONNECT: @data_a 0 0 2 0 data 0 0 2 0
// Retrieval info: CONNECT: @wren_a 0 0 0 0 wren 0 0 0 0
// Retrieval info: CONNECT: q 0 0 2 0 @q_a 0 0 2 0
// Retrieval info: GEN_FILE: TYPE_NORMAL ramTP.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL ramTP.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL ramTP.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL ramTP.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL ramTP_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL ramTP_bb.v TRUE
// Retrieval info: LIB_FILE: altera_mf
