module sequence_recognizer();

endmodule
